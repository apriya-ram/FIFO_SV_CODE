


package fifo_pkg;
//ADD_CODE: `include the fifo_transaction file
  `include "fifo_transaction.sv"
//ADD_CODE: `include the generator.sv file
  `include "generator.sv"
//ADD_CODE: `include the driver.sv file
  `include "driver.sv"
//ADD_CODE: `include the monitor.sv file
  `include "monitor.sv"
//ADD_CODE: `include the scoreboard.sv file
  `include "scoreboard.sv"
//ADD_CODE: `include the environment.sv file
  `include "environment.sv"
//ADD_CODE: `include the test.sv file
  `include "test.sv"
endpackage
